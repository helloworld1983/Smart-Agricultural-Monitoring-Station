----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    17:19:25 03/10/2019 
-- Design Name: 
-- Module Name:    ADC_Input - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use IEEE.NUMERIC_STD;



entity ADC_Input is
  Port		(clk 			: in std_logic;
					 reset 		: in std_logic;
					 switch		: in std_logic;
					 ADC_EN	  : in std_logic;
					 ADC			: in std_logic_vector(7 downto 0);
					 ADC_DONE : out std_logic;
					 ADC_PER  : out std_logic_vector(7 downto 0);
					 ADC_VAL	: out std_logic_vector(31 downto 0);
					 ADC_PER_DISP : out std_logic_vector(31 downto 0));
end ADC_Input;

architecture Behavioral of ADC_Input is

begin
ADC_Lookup:process(clk,reset,switch)

	begin
	if (reset ='1')then
		ADC_VAL<=(others => '0');
		ADC_PER<=(others => '0');
		ADC_PER_DISP<=(others => '0');
		ADC_DONE<='0';
	elsif rising_edge(clk)then
		if(switch='1')then
		 if(ADC_EN='1')then
			case ADC is
				when"00000000"=> ADC_VAL<="10110000001100000101010100000000"; ADC_PER<="00000000"; ADC_PER_DISP<="00110000000000000000000000000000";--0
				when"00000001"=> ADC_VAL<="10110000001100000101010100000000"; ADC_PER<="00000000"; ADC_PER_DISP<="00110000000000000000000000000000";--0.01 
				when"00000010"=> ADC_VAL<="10110000001100000101010100000000"; ADC_PER<="00000000"; ADC_PER_DISP<="00110000000000000000000000000000";--0.02 
				when"00000011"=> ADC_VAL<="10110000001100000101010100000000"; ADC_PER<="00000001"; ADC_PER_DISP<="00110001000000000000000000000000";--0.03 
				when"00000100"=> ADC_VAL<="10110000001100000101010100000000"; ADC_PER<="00000001"; ADC_PER_DISP<="00110001000000000000000000000000";--0.05 
				when"00000101"=> ADC_VAL<="10110000001100000101010100000000"; ADC_PER<="00000001"; ADC_PER_DISP<="00110001000000000000000000000000";--0.06 
				when"00000110"=> ADC_VAL<="10110000001100000101010100000000"; ADC_PER<="00000010"; ADC_PER_DISP<="00110010000000000000000000000000";--0.07 
				when"00000111"=> ADC_VAL<="10110000001100000101010100000000"; ADC_PER<="00000010"; ADC_PER_DISP<="00110010000000000000000000000000";--0.09 
				when"00001000"=> ADC_VAL<="10110000001100010101010100000000"; ADC_PER<="00000011"; ADC_PER_DISP<="00110011000000000000000000000000";--0.10 
				when"00001001"=> ADC_VAL<="10110000001100010101010100000000"; ADC_PER<="00000011"; ADC_PER_DISP<="00110011000000000000000000000000";--0.11 
				when"00001010"=> ADC_VAL<="10110000001100010101010100000000"; ADC_PER<="00000011"; ADC_PER_DISP<="00110011000000000000000000000000";--0.12 
				when"00001011"=> ADC_VAL<="10110000001100010101010100000000"; ADC_PER<="00000100"; ADC_PER_DISP<="00110100000000000000000000000000";--0.14 
				when"00001100"=> ADC_VAL<="10110000001100010101010100000000"; ADC_PER<="00000100"; ADC_PER_DISP<="00110100000000000000000000000000";--0.15 
				when"00001101"=> ADC_VAL<="10110000001100010101010100000000"; ADC_PER<="00000101"; ADC_PER_DISP<="00110101000000000000000000000000";--0.16 
				when"00001110"=> ADC_VAL<="10110000001100010101010100000000"; ADC_PER<="00000101"; ADC_PER_DISP<="00110101000000000000000000000000";--0.18 
				when"00001111"=> ADC_VAL<="10110000001100010101010100000000"; ADC_PER<="00000101"; ADC_PER_DISP<="00110101000000000000000000000000";--0.19 
				when"00010000"=> ADC_VAL<="10110000001100010101010100000000"; ADC_PER<="00000110"; ADC_PER_DISP<="00110110000000000000000000000000";--0.20 
				when"00010001"=> ADC_VAL<="10110000001100010101010100000000"; ADC_PER<="00000110"; ADC_PER_DISP<="00110110000000000000000000000000";--0.22
				when"00010010"=> ADC_VAL<="10110000001100010101010100000000"; ADC_PER<="00000111"; ADC_PER_DISP<="00110111000000000000000000000000";--0.23 
				when"00010011"=> ADC_VAL<="10110000001100010101010100000000"; ADC_PER<="00000111"; ADC_PER_DISP<="00110111000000000000000000000000";--0.24 
				when"00010100"=> ADC_VAL<="10110000001100010101010100000000"; ADC_PER<="00000111"; ADC_PER_DISP<="00110111000000000000000000000000";--0.25 
				when"00010101"=> ADC_VAL<="10110000001100010101010100000000"; ADC_PER<="00001000"; ADC_PER_DISP<="00111000000000000000000000000000";--0.27 
				when"00010110"=> ADC_VAL<="10110000001100010101010100000000"; ADC_PER<="00001000"; ADC_PER_DISP<="00111000000000000000000000000000";--0.28 
				when"00010111"=> ADC_VAL<="10110000001100010101010100000000"; ADC_PER<="00001001"; ADC_PER_DISP<="00111001000000000000000000000000";--0.29 
				when"00011000"=> ADC_VAL<="10110000001100110101010100000000"; ADC_PER<="00001001"; ADC_PER_DISP<="00111001000000000000000000000000";--0.31 
				when"00011001"=> ADC_VAL<="10110000001100110101010100000000"; ADC_PER<="00001001"; ADC_PER_DISP<="00111001000000000000000000000000";--0.32 
				when"00011010"=> ADC_VAL<="10110000001100110101010100000000"; ADC_PER<="00001010"; ADC_PER_DISP<="00110001001100000000000000000000";--0.33 -10%
				when"00011011"=> ADC_VAL<="10110000001100110101010100000000"; ADC_PER<="00001010"; ADC_PER_DISP<="00110001001100000000000000000000";--0.34 
				when"00011100"=> ADC_VAL<="10110000001100110101010100000000"; ADC_PER<="00001010"; ADC_PER_DISP<="00110001001100000000000000000000";--0.36 
				when"00011101"=> ADC_VAL<="10110000001100110101010100000000"; ADC_PER<="00001011"; ADC_PER_DISP<="00110001001100010000000000000000";--0.37 
				when"00011110"=> ADC_VAL<="10110000001100110101010100000000"; ADC_PER<="00001011"; ADC_PER_DISP<="00110001001100010000000000000000";--0.38 
				when"00011111"=> ADC_VAL<="10110000001101000101010100000000"; ADC_PER<="00001100"; ADC_PER_DISP<="00110001001100100000000000000000";--0.40 
				when"00100000"=> ADC_VAL<="10110000001101000101010100000000"; ADC_PER<="00001100"; ADC_PER_DISP<="00110001001100100000000000000000";--0.41 
				when"00100001"=> ADC_VAL<="10110000001101000101010100000000"; ADC_PER<="00001100"; ADC_PER_DISP<="00110001001100100000000000000000";--0.42 
				when"00100010"=> ADC_VAL<="10110000001101000101010100000000"; ADC_PER<="00001101"; ADC_PER_DISP<="00110001001100110000000000000000";--0.44
				when"00100011"=> ADC_VAL<="10110000001101000101010100000000"; ADC_PER<="00001101"; ADC_PER_DISP<="00110001001100110000000000000000";--0.45 
				when"00100100"=> ADC_VAL<="10110000001101000101010100000000"; ADC_PER<="00001110"; ADC_PER_DISP<="00110001001101000000000000000000";--0.46 
				when"00100101"=> ADC_VAL<="10110000001101000101010100000000"; ADC_PER<="00001110"; ADC_PER_DISP<="00110001001101000000000000000000";--0.47 
				when"00100110"=> ADC_VAL<="10110000001101000101010100000000"; ADC_PER<="00001110"; ADC_PER_DISP<="00110001001101000000000000000000";--0.49 
				when"00100111"=> ADC_VAL<="10110000001101010101010100000000"; ADC_PER<="00001111"; ADC_PER_DISP<="00110001001101010000000000000000";--0.50 
				when"00101000"=> ADC_VAL<="10110000001101010101010100000000"; ADC_PER<="00001111"; ADC_PER_DISP<="00110001001101010000000000000000";--0.51 
				when"00101001"=> ADC_VAL<="10110000001101010101010100000000"; ADC_PER<="00010000"; ADC_PER_DISP<="00110001001101100000000000000000";--0.53 
				when"00101010"=> ADC_VAL<="10110000001101010101010100000000"; ADC_PER<="00010000"; ADC_PER_DISP<="00110001001101100000000000000000";--0.54 
				when"00101011"=> ADC_VAL<="10110000001101010101010100000000"; ADC_PER<="00010000"; ADC_PER_DISP<="00110001001101100000000000000000";--0.55 
				when"00101100"=> ADC_VAL<="10110000001101010101010100000000"; ADC_PER<="00010001"; ADC_PER_DISP<="00110001001101110000000000000000";--0.56 
				when"00101101"=> ADC_VAL<="10110000001101010101010100000000"; ADC_PER<="00010001"; ADC_PER_DISP<="00110001001101110000000000000000";--0.58 
				when"00101110"=> ADC_VAL<="10110000001101010101010100000000"; ADC_PER<="00010010"; ADC_PER_DISP<="00110001001110000000000000000000";--0.59 
				when"00101111"=> ADC_VAL<="10110000001101010101010100000000"; ADC_PER<="00010010"; ADC_PER_DISP<="00110001001110000000000000000000";--0.60 
				when"00110000"=> ADC_VAL<="10110000001101010101010100000000"; ADC_PER<="00010010"; ADC_PER_DISP<="00110001001110000000000000000000";--0.62 
				when"00110001"=> ADC_VAL<="10110000001101010101010100000000"; ADC_PER<="00010011"; ADC_PER_DISP<="00110001001110010000000000000000";--0.63 
				when"00110010"=> ADC_VAL<="10110000001101010101010100000000"; ADC_PER<="00010011"; ADC_PER_DISP<="00110001001110010000000000000000";--0.64 
				when"00110011"=> ADC_VAL<="10110000001101010101010100000000"; ADC_PER<="00010100"; ADC_PER_DISP<="00110010001100000000000000000000";--0.66  -20%
				when"00110100"=> ADC_VAL<="10110000001101010101010100000000"; ADC_PER<="00010100"; ADC_PER_DISP<="00110010001100000000000000000000";--0.67 
				when"00110101"=> ADC_VAL<="10110000001101010101010100000000"; ADC_PER<="00010100"; ADC_PER_DISP<="00110010001100000000000000000000";--0.68 
				when"00110110"=> ADC_VAL<="10110000001101010101010100000000"; ADC_PER<="00010101"; ADC_PER_DISP<="00110010001100010000000000000000";--0.69 
				when"00110111"=> ADC_VAL<="10110000001101110101010100000000"; ADC_PER<="00010101"; ADC_PER_DISP<="00110010001100010000000000000000";--0.71 
				when"00111000"=> ADC_VAL<="10110000001101110101010100000000"; ADC_PER<="00010101"; ADC_PER_DISP<="00110010001100010000000000000000";--0.72 
				when"00111001"=> ADC_VAL<="10110000001101110101010100000000"; ADC_PER<="00010110"; ADC_PER_DISP<="00110010001100100000000000000000";--0.73 
				when"00111010"=> ADC_VAL<="10110000001101110101010100000000"; ADC_PER<="00010110"; ADC_PER_DISP<="00110010001100100000000000000000";--0.75 
				when"00111011"=> ADC_VAL<="10110000001101110101010100000000"; ADC_PER<="00010111"; ADC_PER_DISP<="00110010001100110000000000000000";--0.76 
				when"00111100"=> ADC_VAL<="10110000001101110101010100000000"; ADC_PER<="00010111"; ADC_PER_DISP<="00110010001100110000000000000000";--0.77 
				when"00111101"=> ADC_VAL<="10110000001101110101010100000000"; ADC_PER<="00010111"; ADC_PER_DISP<="00110010001100110000000000000000";--0.78 
				when"00111110"=> ADC_VAL<="10110000001110000101010100000000"; ADC_PER<="00011000"; ADC_PER_DISP<="00110010001101000000000000000000";--0.80 
				when"00111111"=> ADC_VAL<="10110000001110000101010100000000"; ADC_PER<="00011000"; ADC_PER_DISP<="00110010001101000000000000000000";--0.81 
				when"01000000"=> ADC_VAL<="10110000001110000101010100000000"; ADC_PER<="00011001"; ADC_PER_DISP<="00110010001101010000000000000000";--0.82 
				when"01000001"=> ADC_VAL<="10110000001110000101010100000000"; ADC_PER<="00011001"; ADC_PER_DISP<="00110010001101010000000000000000";--0.84 
				when"01000010"=> ADC_VAL<="10110000001110000101010100000000"; ADC_PER<="00011001"; ADC_PER_DISP<="00110010001101010000000000000000";--0.85 
				when"01000011"=> ADC_VAL<="10110000001110000101010100000000"; ADC_PER<="00011010"; ADC_PER_DISP<="00110010001101100000000000000000";--0.86 
				when"01000100"=> ADC_VAL<="10110000001110000101010100000000"; ADC_PER<="00011010"; ADC_PER_DISP<="00110010001101100000000000000000";--0.88
				when"01000101"=> ADC_VAL<="10110000001110000101010100000000"; ADC_PER<="00011011"; ADC_PER_DISP<="00110010001101110000000000000000";--0.892941
				when"01000110"=> ADC_VAL<="10110000001110010101010100000000"; ADC_PER<="00011011"; ADC_PER_DISP<="00110010001101110000000000000000";--0.905883
				when"01000111"=> ADC_VAL<="10110000001110010101010100000000"; ADC_PER<="00011011"; ADC_PER_DISP<="00110010001101110000000000000000";--0.918824
				when"01001000"=> ADC_VAL<="10110000001110010101010100000000"; ADC_PER<="00011100"; ADC_PER_DISP<="00110010001110000000000000000000";--0.931765
				when"01001001"=> ADC_VAL<="10110000001110010101010100000000"; ADC_PER<="00011100"; ADC_PER_DISP<="00110010001110000000000000000000";--0.944706
				when"01001010"=> ADC_VAL<="10110000001110010101010100000000"; ADC_PER<="00011101"; ADC_PER_DISP<="00110010001110010000000000000000";--0.957647
				when"01001011"=> ADC_VAL<="10110000001110010101010100000000"; ADC_PER<="00011101"; ADC_PER_DISP<="00110010001110010000000000000000";--0.970589
				when"01001100"=> ADC_VAL<="10110000001110010101010100000000"; ADC_PER<="00011101"; ADC_PER_DISP<="00110010001110010000000000000000";--0.98353
				when"01001101"=> ADC_VAL<="10110000001110010101010100000000"; ADC_PER<="00011110"; ADC_PER_DISP<="00110011001100000000000000000000";--0.996471 --30%
				when"01001110"=> ADC_VAL<="10110001001100000101010100000000"; ADC_PER<="00011110"; ADC_PER_DISP<="00110011001100000000000000000000";--1.00941
				when"01001111"=> ADC_VAL<="10110001001100000101010100000000"; ADC_PER<="00011110"; ADC_PER_DISP<="00110011001100000000000000000000";--1.02235
				when"01010000"=> ADC_VAL<="10110001001100000101010100000000"; ADC_PER<="00011111"; ADC_PER_DISP<="00110011001100010000000000000000";--1.03529
				when"01010001"=> ADC_VAL<="10110001001100000101010100000000"; ADC_PER<="00011111"; ADC_PER_DISP<="00110011001100010000000000000000";--1.04824
				when"01010010"=> ADC_VAL<="10110001001100000101010100000000"; ADC_PER<="00100000"; ADC_PER_DISP<="00110011001100100000000000000000";--1.06118
				when"01010011"=> ADC_VAL<="10110001001100000101010100000000"; ADC_PER<="00100000"; ADC_PER_DISP<="00110011001100100000000000000000";--1.07412
				when"01010100"=> ADC_VAL<="10110001001100000101010100000000"; ADC_PER<="00100000"; ADC_PER_DISP<="00110011001100100000000000000000";--1.08706
				when"01010101"=> ADC_VAL<="10110001001100010101010100000000"; ADC_PER<="00100001"; ADC_PER_DISP<="00110011001100110000000000000000";--1.1
				when"01010110"=> ADC_VAL<="10110001001100010101010100000000"; ADC_PER<="00100001"; ADC_PER_DISP<="00110011001100110000000000000000";--1.11294
				when"01010111"=> ADC_VAL<="10110001001100010101010100000000"; ADC_PER<="00100010"; ADC_PER_DISP<="00110011001101000000000000000000";--1.12588
				when"01011000"=> ADC_VAL<="10110001001100010101010100000000"; ADC_PER<="00100010"; ADC_PER_DISP<="00110011001101000000000000000000";--1.13882
				when"01011001"=> ADC_VAL<="10110001001100010101010100000000"; ADC_PER<="00100010"; ADC_PER_DISP<="00110011001101000000000000000000";--1.15176
				when"01011010"=> ADC_VAL<="10110001001100010101010100000000"; ADC_PER<="00100011"; ADC_PER_DISP<="00110011001101010000000000000000";--1.16471
				when"01011011"=> ADC_VAL<="10110001001100010101010100000000"; ADC_PER<="00100011"; ADC_PER_DISP<="00110011001101010000000000000000";--1.17765
				when"01011100"=> ADC_VAL<="10110001001100010101010100000000"; ADC_PER<="00100100"; ADC_PER_DISP<="00110011001101100000000000000000";--1.19059
				when"01011101"=> ADC_VAL<="10110001001100010101010100000000"; ADC_PER<="00100100"; ADC_PER_DISP<="00110011001101100000000000000000";--1.20353
				when"01011110"=> ADC_VAL<="10110001001100010101010100000000"; ADC_PER<="00100100"; ADC_PER_DISP<="00110011001101100000000000000000";--1.21647
				when"01011111"=> ADC_VAL<="10110001001100010101010100000000"; ADC_PER<="00100101"; ADC_PER_DISP<="00110011001101110000000000000000";--1.22941
				when"01100000"=> ADC_VAL<="10110001001100010101010100000000"; ADC_PER<="00100101"; ADC_PER_DISP<="00110011001101110000000000000000";--1.24235
				when"01100001"=> ADC_VAL<="10110001001100010101010100000000"; ADC_PER<="00100110"; ADC_PER_DISP<="00110011001110000000000000000000";--1.25529
				when"01100010"=> ADC_VAL<="10110001001100010101010100000000"; ADC_PER<="00100110"; ADC_PER_DISP<="00110011001110000000000000000000";--1.26823
				when"01100011"=> ADC_VAL<="10110001001100010101010100000000"; ADC_PER<="00100110"; ADC_PER_DISP<="00110011001110000000000000000000";--1.28118
				when"01100100"=> ADC_VAL<="10110001001100010101010100000000"; ADC_PER<="00100111"; ADC_PER_DISP<="00110011001110010000000000000000";--1.29412
				when"01100101"=> ADC_VAL<="10110001001100110101010100000000"; ADC_PER<="00100111"; ADC_PER_DISP<="00110011001110010000000000000000";--1.30706
				when"01100110"=> ADC_VAL<="10110001001100110101010100000000"; ADC_PER<="00101000"; ADC_PER_DISP<="00110100001100000000000000000000";--1.32    --40%
				when"01100111"=> ADC_VAL<="10110001001100110101010100000000"; ADC_PER<="00101000"; ADC_PER_DISP<="00110100001100000000000000000000";--1.33294
				when"01101000"=> ADC_VAL<="10110001001100110101010100000000"; ADC_PER<="00101000"; ADC_PER_DISP<="00110100001100000000000000000000";--1.34588
				when"01101001"=> ADC_VAL<="10110001001100110101010100000000"; ADC_PER<="00101001"; ADC_PER_DISP<="00110100001100010000000000000000";--1.35882
				when"01101010"=> ADC_VAL<="10110001001100110101010100000000"; ADC_PER<="00101001"; ADC_PER_DISP<="00110100001100010000000000000000";--1.37176
				when"01101011"=> ADC_VAL<="10110001001100110101010100000000"; ADC_PER<="00101001"; ADC_PER_DISP<="00110100001100010000000000000000";--1.3847
				when"01101100"=> ADC_VAL<="10110001001100110101010100000000"; ADC_PER<="00101010"; ADC_PER_DISP<="00110100001100100000000000000000";--1.39765
				when"01101101"=> ADC_VAL<="10110001001101000101010100000000"; ADC_PER<="00101010"; ADC_PER_DISP<="00110100001100100000000000000000";--1.41059
				when"01101110"=> ADC_VAL<="10110001001101000101010100000000"; ADC_PER<="00101011"; ADC_PER_DISP<="00110100001100110000000000000000";--1.42353
				when"01101111"=> ADC_VAL<="10110001001101000101010100000000"; ADC_PER<="00101011"; ADC_PER_DISP<="00110100001100110000000000000000";--1.43647
				when"01110000"=> ADC_VAL<="10110001001101000101010100000000"; ADC_PER<="00101011"; ADC_PER_DISP<="00110100001100110000000000000000";--1.44941
				when"01110001"=> ADC_VAL<="10110001001101000101010100000000"; ADC_PER<="00101100"; ADC_PER_DISP<="00110100001101000000000000000000";--1.46235
				when"01110010"=> ADC_VAL<="10110001001101000101010100000000"; ADC_PER<="00101100"; ADC_PER_DISP<="00110100001101000000000000000000";--1.47529
				when"01110011"=> ADC_VAL<="10110001001101000101010100000000"; ADC_PER<="00101101"; ADC_PER_DISP<="00110100001101010000000000000000";--1.48823
				when"01110100"=> ADC_VAL<="10110001001101010101010100000000"; ADC_PER<="00101101"; ADC_PER_DISP<="00110100001101010000000000000000";--1.50117
				when"01110101"=> ADC_VAL<="10110001001101010101010100000000"; ADC_PER<="00101101"; ADC_PER_DISP<="00110100001101010000000000000000";--1.51412
				when"01110110"=> ADC_VAL<="10110001001101010101010100000000"; ADC_PER<="00101110"; ADC_PER_DISP<="00110100001101100000000000000000";--1.52706
				when"01110111"=> ADC_VAL<="10110001001101010101010100000000"; ADC_PER<="00101110"; ADC_PER_DISP<="00110100001101100000000000000000";--1.54
				when"01111000"=> ADC_VAL<="10110001001101010101010100000000"; ADC_PER<="00101111"; ADC_PER_DISP<="00110100001101110000000000000000";--1.55294
				when"01111001"=> ADC_VAL<="10110001001101010101010100000000"; ADC_PER<="00101111"; ADC_PER_DISP<="00110100001101110000000000000000";--1.56588
				when"01111010"=> ADC_VAL<="10110001001101010101010100000000"; ADC_PER<="00101111"; ADC_PER_DISP<="00110100001101110000000000000000";--1.57882
				when"01111011"=> ADC_VAL<="10110001001101010101010100000000"; ADC_PER<="00110000"; ADC_PER_DISP<="00110100001110000000000000000000";--1.59176
				when"01111100"=> ADC_VAL<="10110001001101010101010100000000"; ADC_PER<="00110000"; ADC_PER_DISP<="00110100001110000000000000000000";--1.6047
				when"01111101"=> ADC_VAL<="10110001001101010101010100000000"; ADC_PER<="00110001"; ADC_PER_DISP<="00110100001110010000000000000000";--1.61764
				when"01111110"=> ADC_VAL<="10110001001101010101010100000000"; ADC_PER<="00110001"; ADC_PER_DISP<="00110100001110010000000000000000";--1.63059
				when"01111111"=> ADC_VAL<="10110001001101010101010100000000"; ADC_PER<="00110001"; ADC_PER_DISP<="00110100001110010000000000000000";--1.64353
				when"10000000"=> ADC_VAL<="10110001001101010101010100000000"; ADC_PER<="00110010"; ADC_PER_DISP<="00110101001100000000000000000000";--1.65647 --50%
				when"10000001"=> ADC_VAL<="10110001001101010101010100000000"; ADC_PER<="00110010"; ADC_PER_DISP<="00110101001100000000000000000000";--1.66941
				when"10000010"=> ADC_VAL<="10110001001101010101010100000000"; ADC_PER<="00110010"; ADC_PER_DISP<="00110101001100000000000000000000";--1.68235
				when"10000011"=> ADC_VAL<="10110001001101010101010100000000"; ADC_PER<="00110011"; ADC_PER_DISP<="00110101001100010000000000000000";--1.69529
				when"10000100"=> ADC_VAL<="10110001001101110101010100000000"; ADC_PER<="00110011"; ADC_PER_DISP<="00110101001100010000000000000000";---1.70823
				when"10000101"=> ADC_VAL<="10110001001101110101010100000000"; ADC_PER<="00110100"; ADC_PER_DISP<="00110101001100100000000000000000";--1.72117
				when"10000110"=> ADC_VAL<="10110001001101110101010100000000"; ADC_PER<="00110100"; ADC_PER_DISP<="00110101001100100000000000000000";--1.73411
				when"10000111"=> ADC_VAL<="10110001001101110101010100000000"; ADC_PER<="00110100"; ADC_PER_DISP<="00110101001100100000000000000000";--1.74706
				when"10001000"=> ADC_VAL<="10110001001101110101010100000000"; ADC_PER<="00110101"; ADC_PER_DISP<="00110101001100110000000000000000";--1.76
				when"10001001"=> ADC_VAL<="10110001001101110101010100000000"; ADC_PER<="00110101"; ADC_PER_DISP<="00110101001100110000000000000000";--1.77294
				when"10001010"=> ADC_VAL<="10110001001101110101010100000000"; ADC_PER<="00110110"; ADC_PER_DISP<="00110101001101000000000000000000";--1.78588
				when"10001011"=> ADC_VAL<="10110001001101110101010100000000"; ADC_PER<="00110110"; ADC_PER_DISP<="00110101001101000000000000000000";--1.79882
				when"10001100"=> ADC_VAL<="10110001001110000101010100000000"; ADC_PER<="00110110"; ADC_PER_DISP<="00110101001101000000000000000000";--1.81176
				when"10001101"=> ADC_VAL<="10110001001110000101010100000000"; ADC_PER<="00110111"; ADC_PER_DISP<="00110101001101010000000000000000";--1.8247
				when"10001110"=> ADC_VAL<="10110001001110000101010100000000"; ADC_PER<="00110111"; ADC_PER_DISP<="00110101001101010000000000000000";--1.83764
				when"10001111"=> ADC_VAL<="10110001001110000101010100000000"; ADC_PER<="00111000"; ADC_PER_DISP<="00110101001101100000000000000000";--1.85058
				when"10010000"=> ADC_VAL<="10110001001110000101010100000000"; ADC_PER<="00111000"; ADC_PER_DISP<="00110101001101100000000000000000";--1.86353
				when"10010001"=> ADC_VAL<="10110001001110000101010100000000"; ADC_PER<="00111000"; ADC_PER_DISP<="00110101001101100000000000000000";--1.87647
				when"10010010"=> ADC_VAL<="10110001001110000101010100000000"; ADC_PER<="00111001"; ADC_PER_DISP<="00110101001101110000000000000000";--1.88941
				when"10010011"=> ADC_VAL<="10110001001110010101010100000000"; ADC_PER<="00111001"; ADC_PER_DISP<="00110101001101110000000000000000";--1.90235
				when"10010100"=> ADC_VAL<="10110001001110010101010100000000"; ADC_PER<="00111010"; ADC_PER_DISP<="00110101001110000000000000000000";--1.91529
				when"10010101"=> ADC_VAL<="10110001001110010101010100000000"; ADC_PER<="00111010"; ADC_PER_DISP<="00110101001110000000000000000000";--1.92823
				when"10010110"=> ADC_VAL<="10110001001110010101010100000000"; ADC_PER<="00111010"; ADC_PER_DISP<="00110101001110000000000000000000";--1.94117
				when"10010111"=> ADC_VAL<="10110001001110010101010100000000"; ADC_PER<="00111011"; ADC_PER_DISP<="00110101001110010000000000000000";--1.95411
				when"10011000"=> ADC_VAL<="10110001001110010101010100000000"; ADC_PER<="00111011"; ADC_PER_DISP<="00110101001110010000000000000000";--1.96706 
				when"10011001"=> ADC_VAL<="10110001001110010101010100000000"; ADC_PER<="00111100"; ADC_PER_DISP<="00110110001100000000000000000000";--1.98    --60%
				when"10011010"=> ADC_VAL<="10110001001110010101010100000000"; ADC_PER<="00111100"; ADC_PER_DISP<="00110110001100000000000000000000";--1.99294
				when"10011011"=> ADC_VAL<="10110010001100000101010100000000"; ADC_PER<="00111100"; ADC_PER_DISP<="00110110001100000000000000000000";--2.00588
				when"10011100"=> ADC_VAL<="10110010001100000101010100000000"; ADC_PER<="00111101"; ADC_PER_DISP<="00110110001100010000000000000000";--2.01882
				when"10011101"=> ADC_VAL<="10110010001100000101010100000000"; ADC_PER<="00111101"; ADC_PER_DISP<="00110110001100010000000000000000";--2.03176
				when"10011110"=> ADC_VAL<="10110010001100000101010100000000"; ADC_PER<="00111101"; ADC_PER_DISP<="00110110001100010000000000000000";--2.0447
				when"10011111"=> ADC_VAL<="10110010001100000101010100000000"; ADC_PER<="00111110"; ADC_PER_DISP<="00110110001100100000000000000000";--2.05764
				when"10100000"=> ADC_VAL<="10110010001100000101010100000000"; ADC_PER<="00111110"; ADC_PER_DISP<="00110110001100100000000000000000";--2.07058
				when"10100001"=> ADC_VAL<="10110010001100000101010100000000"; ADC_PER<="00111111"; ADC_PER_DISP<="00110110001100110000000000000000";--2.08353
				when"10100010"=> ADC_VAL<="10110010001100000101010100000000"; ADC_PER<="00111111"; ADC_PER_DISP<="00110110001100110000000000000000";--2.09647
				when"10100011"=> ADC_VAL<="10110010001100010101010100000000"; ADC_PER<="00111111"; ADC_PER_DISP<="00110110001100110000000000000000";--2.10941
				when"10100100"=> ADC_VAL<="10110010001100010101010100000000"; ADC_PER<="01000000"; ADC_PER_DISP<="00110110001101000000000000000000";--2.12235
				when"10100101"=> ADC_VAL<="10110010001100010101010100000000"; ADC_PER<="01000000"; ADC_PER_DISP<="00110110001101000000000000000000";--2.13529
				when"10100110"=> ADC_VAL<="10110010001100010101010100000000"; ADC_PER<="01000001"; ADC_PER_DISP<="00110110001101010000000000000000";--2.14823
				when"10100111"=> ADC_VAL<="10110010001100010101010100000000"; ADC_PER<="01000001"; ADC_PER_DISP<="00110110001101010000000000000000";--2.16117
				when"10101000"=> ADC_VAL<="10110010001100010101010100000000"; ADC_PER<="01000001"; ADC_PER_DISP<="00110110001101010000000000000000";--2.17411
				when"10101001"=> ADC_VAL<="10110010001100010101010100000000"; ADC_PER<="01000010"; ADC_PER_DISP<="00110110001101100000000000000000";--2.18705
				when"10101010"=> ADC_VAL<="10110010001100010101010100000000"; ADC_PER<="01000010"; ADC_PER_DISP<="00110110001101100000000000000000";--2.2
				when"10101011"=> ADC_VAL<="10110010001100010101010100000000"; ADC_PER<="01000011"; ADC_PER_DISP<="00110110001101110000000000000000";--2.21294
				when"10101100"=> ADC_VAL<="10110010001100010101010100000000"; ADC_PER<="01000011"; ADC_PER_DISP<="00110110001101110000000000000000";--2.22588
				when"10101101"=> ADC_VAL<="10110010001100010101010100000000"; ADC_PER<="01000011"; ADC_PER_DISP<="00110110001101110000000000000000";--2.23882
				when"10101110"=> ADC_VAL<="10110010001100010101010100000000"; ADC_PER<="01000100"; ADC_PER_DISP<="00110110001110000000000000000000";--2.25176
				when"10101111"=> ADC_VAL<="10110010001100010101010100000000"; ADC_PER<="01000100"; ADC_PER_DISP<="00110110001110000000000000000000";--2.2647
				when"10110000"=> ADC_VAL<="10110010001100010101010100000000"; ADC_PER<="01000101"; ADC_PER_DISP<="00110110001110010000000000000000";--2.27764
				when"10110001"=> ADC_VAL<="10110010001100010101010100000000"; ADC_PER<="01000101"; ADC_PER_DISP<="00110110001110010000000000000000";--2.29058
				when"10110010"=> ADC_VAL<="10110010001100110101010100000000"; ADC_PER<="01000101"; ADC_PER_DISP<="00110110001110010000000000000000";--2.30352
				when"10110011"=> ADC_VAL<="10110010001100110101010100000000"; ADC_PER<="01000110"; ADC_PER_DISP<="00110111001100000000000000000000";--2.31647 --70%
				when"10110100"=> ADC_VAL<="10110010001100110101010100000000"; ADC_PER<="01000110"; ADC_PER_DISP<="00110111001100000000000000000000";--2.32941
				when"10110101"=> ADC_VAL<="10110010001100110101010100000000"; ADC_PER<="01000110"; ADC_PER_DISP<="00110111001100000000000000000000";--2.34235
				when"10110110"=> ADC_VAL<="10110010001100110101010100000000"; ADC_PER<="01000111"; ADC_PER_DISP<="00110111001100010000000000000000";--2.35529
				when"10110111"=> ADC_VAL<="10110010001100110101010100000000"; ADC_PER<="01000111"; ADC_PER_DISP<="00110111001100010000000000000000";--2.36823
				when"10111000"=> ADC_VAL<="10110010001100110101010100000000"; ADC_PER<="01001000"; ADC_PER_DISP<="00110111001100100000000000000000";--2.38117
				when"10111001"=> ADC_VAL<="10110010001100110101010100000000"; ADC_PER<="01001000"; ADC_PER_DISP<="00110111001100100000000000000000";--2.39411
				when"10111010"=> ADC_VAL<="10110010001101000101010100000000"; ADC_PER<="01001000"; ADC_PER_DISP<="00110111001100100000000000000000";--2.40705
				when"10111011"=> ADC_VAL<="10110010001101000101010100000000"; ADC_PER<="01001001"; ADC_PER_DISP<="00110111001100110000000000000000";--2.41999
				when"10111100"=> ADC_VAL<="10110010001101000101010100000000"; ADC_PER<="01001001"; ADC_PER_DISP<="00110111001100110000000000000000";--2.43294
				when"10111101"=> ADC_VAL<="10110010001101000101010100000000"; ADC_PER<="01001010"; ADC_PER_DISP<="00110111001101000000000000000000";--2.44588
				when"10111110"=> ADC_VAL<="10110010001101000101010100000000"; ADC_PER<="01001010"; ADC_PER_DISP<="00110111001101000000000000000000";--2.45882
				when"10111111"=> ADC_VAL<="10110010001101000101010100000000"; ADC_PER<="01001010"; ADC_PER_DISP<="00110111001101000000000000000000";--2.47176
				when"11000000"=> ADC_VAL<="10110010001101000101010100000000"; ADC_PER<="01001011"; ADC_PER_DISP<="00110111001101010000000000000000";--2.4847
				when"11000001"=> ADC_VAL<="10110010001101000101010100000000"; ADC_PER<="01001011"; ADC_PER_DISP<="00110111001101010000000000000000";--2.49764
				when"11000010"=> ADC_VAL<="10110010001101010101010100000000"; ADC_PER<="01001100"; ADC_PER_DISP<="00110111001101100000000000000000";--2.51058
				when"11000011"=> ADC_VAL<="10110010001101010101010100000000"; ADC_PER<="01001100"; ADC_PER_DISP<="00110111001101100000000000000000";--2.52352
				when"11000100"=> ADC_VAL<="10110010001101010101010100000000"; ADC_PER<="01001100"; ADC_PER_DISP<="00110111001101100000000000000000";--2.53646
				when"11000101"=> ADC_VAL<="10110010001101010101010100000000"; ADC_PER<="01001101"; ADC_PER_DISP<="00110111001101110000000000000000";--2.54941
				when"11000110"=> ADC_VAL<="10110010001101010101010100000000"; ADC_PER<="01001101"; ADC_PER_DISP<="00110111001101110000000000000000";--2.56235
				when"11000111"=> ADC_VAL<="10110010001101010101010100000000"; ADC_PER<="01001110"; ADC_PER_DISP<="00110111001110000000000000000000";--2.57529
				when"11001000"=> ADC_VAL<="10110010001101010101010100000000"; ADC_PER<="01001110"; ADC_PER_DISP<="00110111001110000000000000000000";--2.58823
				when"11001001"=> ADC_VAL<="10110010001101010101010100000000"; ADC_PER<="01001110"; ADC_PER_DISP<="00110111001110000000000000000000";--2.60117
				when"11001010"=> ADC_VAL<="10110010001101010101010100000000"; ADC_PER<="01001111"; ADC_PER_DISP<="00110111001110010000000000000000";--2.61411
				when"11001011"=> ADC_VAL<="10110010001101010101010100000000"; ADC_PER<="01001111"; ADC_PER_DISP<="00110111001110010000000000000000";--2.62705
				when"11001100"=> ADC_VAL<="10110010001101010101010100000000"; ADC_PER<="01010000"; ADC_PER_DISP<="00111000001100000000000000000000";--2.63999 --80%
				when"11001101"=> ADC_VAL<="10110010001101010101010100000000"; ADC_PER<="01010000"; ADC_PER_DISP<="00111000001100000000000000000000";--2.65293
				when"11001110"=> ADC_VAL<="10110010001101010101010100000000"; ADC_PER<="01010000"; ADC_PER_DISP<="00111000001100000000000000000000";--2.66588
				when"11001111"=> ADC_VAL<="10110010001101010101010100000000"; ADC_PER<="01010001"; ADC_PER_DISP<="00111000001100010000000000000000";--2.67882
				when"11010000"=> ADC_VAL<="10110010001101010101010100000000"; ADC_PER<="01010001"; ADC_PER_DISP<="00111000001100010000000000000000";--2.69176
				when"11010001"=> ADC_VAL<="10110010001101110101010100000000"; ADC_PER<="01010001"; ADC_PER_DISP<="00111000001100010000000000000000";--2.7047
				when"11010010"=> ADC_VAL<="10110010001101110101010100000000"; ADC_PER<="01010010"; ADC_PER_DISP<="00111000001100100000000000000000";--2.71764
				when"11010011"=> ADC_VAL<="10110010001101110101010100000000"; ADC_PER<="01010010"; ADC_PER_DISP<="00111000001100100000000000000000";--2.73058
				when"11010100"=> ADC_VAL<="10110010001101110101010100000000"; ADC_PER<="01010011"; ADC_PER_DISP<="00111000001100110000000000000000";--2.74352
				when"11010101"=> ADC_VAL<="10110010001101110101010100000000"; ADC_PER<="01010011"; ADC_PER_DISP<="00111000001100110000000000000000";--2.75646
				when"11010110"=> ADC_VAL<="10110010001101110101010100000000"; ADC_PER<="01010011"; ADC_PER_DISP<="00111000001100110000000000000000";--2.7694
				when"11010111"=> ADC_VAL<="10110010001101110101010100000000"; ADC_PER<="01010100"; ADC_PER_DISP<="00111000001101000000000000000000";--2.78235
				when"11011000"=> ADC_VAL<="10110010001101110101010100000000"; ADC_PER<="01010100"; ADC_PER_DISP<="00111000001101000000000000000000";--2.79529
				when"11011001"=> ADC_VAL<="10110010001110000101010100000000"; ADC_PER<="01010101"; ADC_PER_DISP<="00111000001101010000000000000000";--2.80823
				when"11011010"=> ADC_VAL<="10110010001110000101010100000000"; ADC_PER<="01010101"; ADC_PER_DISP<="00111000001101010000000000000000";--2.82117
				when"11011011"=> ADC_VAL<="10110010001110000101010100000000"; ADC_PER<="01010101"; ADC_PER_DISP<="00111000001101010000000000000000";--2.83411
				when"11011100"=> ADC_VAL<="10110010001110000101010100000000"; ADC_PER<="01010110"; ADC_PER_DISP<="00111000001101100000000000000000";--2.84705
				when"11011101"=> ADC_VAL<="10110010001110000101010100000000"; ADC_PER<="01010110"; ADC_PER_DISP<="00111000001101100000000000000000";--2.85999
				when"11011110"=> ADC_VAL<="10110010001110000101010100000000"; ADC_PER<="01010111"; ADC_PER_DISP<="00111000001101110000000000000000";--2.87293
				when"11011111"=> ADC_VAL<="10110010001110000101010100000000"; ADC_PER<="01010111"; ADC_PER_DISP<="00111000001101110000000000000000";--2.88587
				when"11100000"=> ADC_VAL<="10110010001110000101010100000000"; ADC_PER<="01010111"; ADC_PER_DISP<="00111000001101110000000000000000";--2.89882
				when"11100001"=> ADC_VAL<="10110010001110010101010100000000"; ADC_PER<="01011000"; ADC_PER_DISP<="00111000001110000000000000000000";--2.91176
				when"11100010"=> ADC_VAL<="10110010001110010101010100000000"; ADC_PER<="01011000"; ADC_PER_DISP<="00111000001110000000000000000000";--2.9247
				when"11100011"=> ADC_VAL<="10110010001110010101010100000000"; ADC_PER<="01011001"; ADC_PER_DISP<="00111000001110010000000000000000";--2.93764
				when"11100100"=> ADC_VAL<="10110010001110010101010100000000"; ADC_PER<="01011001"; ADC_PER_DISP<="00111000001110010000000000000000";--2.95058
				when"11100101"=> ADC_VAL<="10110010001110010101010100000000"; ADC_PER<="01011001"; ADC_PER_DISP<="00111000001110010000000000000000";--2.96352
				when"11100110"=> ADC_VAL<="10110010001110010101010100000000"; ADC_PER<="01011010"; ADC_PER_DISP<="00111001001100000000000000000000";--2.97646 --90%
				when"11100111"=> ADC_VAL<="10110010001110010101010100000000"; ADC_PER<="01011010"; ADC_PER_DISP<="00111001001100000000000000000000";--2.9894
				when"11101000"=> ADC_VAL<="10110011001100000101010100000000"; ADC_PER<="01011010"; ADC_PER_DISP<="00111001001100000000000000000000";--3.00234
				when"11101001"=> ADC_VAL<="10110011001100000101010100000000"; ADC_PER<="01011011"; ADC_PER_DISP<="00111001001100010000000000000000";--3.01529
				when"11101010"=> ADC_VAL<="10110011001100000101010100000000"; ADC_PER<="01011011"; ADC_PER_DISP<="00111001001100010000000000000000";--3.02823
				when"11101011"=> ADC_VAL<="10110011001100000101010100000000"; ADC_PER<="01011100"; ADC_PER_DISP<="00111001001100100000000000000000";--3.04117
				when"11101100"=> ADC_VAL<="10110011001100000101010100000000"; ADC_PER<="01011100"; ADC_PER_DISP<="00111001001100100000000000000000";--3.05411
				when"11101101"=> ADC_VAL<="10110011001100000101010100000000"; ADC_PER<="01011100"; ADC_PER_DISP<="00111001001100100000000000000000";--3.06705
				when"11101110"=> ADC_VAL<="10110011001100000101010100000000"; ADC_PER<="01011101"; ADC_PER_DISP<="00111001001100110000000000000000";--3.07999
				when"11101111"=> ADC_VAL<="10110011001100000101010100000000"; ADC_PER<="01011101"; ADC_PER_DISP<="00111001001100110000000000000000";--3.09293
				when"11110000"=> ADC_VAL<="10110011001100010101010100000000"; ADC_PER<="01011110"; ADC_PER_DISP<="00111001001101000000000000000000";--3.10587
				when"11110001"=> ADC_VAL<="10110011001100010101010100000000"; ADC_PER<="01011110"; ADC_PER_DISP<="00111001001101000000000000000000";--3.11881
				when"11110010"=> ADC_VAL<="10110011001100010101010100000000"; ADC_PER<="01011110"; ADC_PER_DISP<="00111001001101000000000000000000";--3.13176
				when"11110011"=> ADC_VAL<="10110011001100010101010100000000"; ADC_PER<="01011111"; ADC_PER_DISP<="00111001001101010000000000000000";--3.1447
				when"11110100"=> ADC_VAL<="10110011001100010101010100000000"; ADC_PER<="01011111"; ADC_PER_DISP<="00111001001101010000000000000000";--3.15764
				when"11110101"=> ADC_VAL<="10110011001100010101010100000000"; ADC_PER<="01100000"; ADC_PER_DISP<="00111001001101100000000000000000";--3.17058
				when"11110110"=> ADC_VAL<="10110011001100010101010100000000"; ADC_PER<="01100000"; ADC_PER_DISP<="00111001001101100000000000000000";--3.18352
				when"11110111"=> ADC_VAL<="10110011001100010101010100000000"; ADC_PER<="01100000"; ADC_PER_DISP<="00111001001101100000000000000000";--3.19646
				when"11111000"=> ADC_VAL<="10110011001100010101010100000000"; ADC_PER<="01100001"; ADC_PER_DISP<="00111001001101110000000000000000";--3.2094
				when"11111001"=> ADC_VAL<="10110011001100010101010100000000"; ADC_PER<="01100001"; ADC_PER_DISP<="00111001001101110000000000000000";--3.22234
				when"11111010"=> ADC_VAL<="10110011001100010101010100000000"; ADC_PER<="01100010"; ADC_PER_DISP<="00111001001110000000000000000000";--3.23529
				when"11111011"=> ADC_VAL<="10110011001100010101010100000000"; ADC_PER<="01100010"; ADC_PER_DISP<="00111001001110000000000000000000";--3.24823
				when"11111100"=> ADC_VAL<="10110011001100010101010100000000"; ADC_PER<="01100010"; ADC_PER_DISP<="00111001001110000000000000000000";--3.26117
				when"11111101"=> ADC_VAL<="10110011001100010101010100000000"; ADC_PER<="01100011"; ADC_PER_DISP<="00111001001110010000000000000000";--3.27411
				when"11111110"=> ADC_VAL<="10110011001100010101010100000000"; ADC_PER<="01100011"; ADC_PER_DISP<="00111001001110010000000000000000";--3.28705
				when"11111111"=> ADC_VAL<="10110011001100010101010100000000"; ADC_PER<="01100100"; ADC_PER_DISP<="00111001001110010000000000000000";--3.29999
				when others =>ADC_VAL<= (others => '0'); ADC_PER<= (others => '0');
			end case;
			ADC_DONE<='1';
		 elsif(ADC_EN='0')then
			ADC_DONE<='0';
		 end if;
		end if;
	end if;
end process;
	
	
end Behavioral;

